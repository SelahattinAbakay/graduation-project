`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.01.2024 23:08:45
// Design Name: 
// Module Name: DECODE
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module decode_cycle(
input        clk,
input [7:0]  address_from_data_out_ff,
output [7:0] result_rdA,result_rdB
);
wire [7:0] rdA,rdB;
DECODE decoder_module(.clk(clk),.address_from_data_out_ff(address_from_data_out_ff),.rdA(rdA),.rdB(rdB));
mux_rdA multiplexerrdA(.rdA(rdA),.result_rdA(result_rdA));
mux_rdB multiplexerrdB(.rdB(rdB),.result_rdB(result_rdB));
endmodule

module DECODE(
input clk,
input [7:0] address_from_data_out_ff,
output reg [7:0] rdA,
output reg [7:0] rdB
    );   
always@(posedge clk)
begin
case(address_from_data_out_ff)
8'b00000000: rdA <= 8'b00000000  ;
8'b00000001: rdA <= 8'b00000001  ;
8'b00000010: rdA <= 8'b00000010  ;
8'b00000011: rdA <= 8'b00000011  ;
8'b00000100: rdA <= 8'b00000100  ;
8'b00000101: rdA <= 8'b00000101  ;
8'b00000110: rdA <= 8'b00000110  ;
8'b00000111: rdA <= 8'b00000111  ;
8'b00001000: rdA <= 8'b00001000  ;
8'b00001001: rdA <= 8'b00001001  ;
8'b00001010: rdA <= 8'b00001010  ;
8'b00001011: rdA <= 8'b00001011  ;
8'b00001100: rdA <= 8'b00001100  ;
8'b00001101: rdA <= 8'b00001101  ;
8'b00001110: rdA <= 8'b00001110  ;
8'b00001111: rdA <= 8'b00001111  ;
8'b00010000: rdA <= 8'b00010000;
8'b00010001: rdA <= 8'b00010001;
8'b00010010: rdA <= 8'b00010010;
8'b00010011: rdA <= 8'b00010011;
8'b00010100: rdA <= 8'b00010100;
8'b00010101: rdA <= 8'b00010101;
8'b00010110: rdA <= 8'b00010110;
8'b00010111: rdA <= 8'b00010111;
8'b00011000: rdA <= 8'b00011000;
8'b00011001: rdA <= 8'b00011001;
8'b00011010: rdA <= 8'b00011010;
8'b00011011: rdA <= 8'b00011011;
8'b00011100: rdA <= 8'b00011100;
8'b00011101: rdA <= 8'b00011101;
8'b00011110: rdA <= 8'b00011110;
8'b00011111: rdA <= 8'b00011111;
8'b00100000: rdA <= 8'b00100000;
8'b00100001: rdA <= 8'b00100001;
8'b00100010: rdA <= 8'b00100010;
8'b00100011: rdA <= 8'b00100011;
8'b00100100: rdA <= 8'b00100100;
8'b00100101: rdA <= 8'b00100101;
8'b00100110: rdA <= 8'b00100110;
8'b00100111: rdA <= 8'b00100111;
8'b00101000: rdA <= 8'b00101000;
8'b00101001: rdA <= 8'b00101001;
8'b00101010: rdA <= 8'b00101010;
8'b00101011: rdA <= 8'b00101011;
8'b00101100: rdA <= 8'b00101100;
8'b00101101: rdA <= 8'b00101101;
8'b00101110: rdA <= 8'b00101110;
8'b00101111: rdA <= 8'b00101111;
8'b00110000: rdA <= 8'b00110000;
8'b00110001: rdA <= 8'b00110001;
8'b00110010: rdA <= 8'b00110010;
8'b00110011: rdA <= 8'b00110011;
8'b00110100: rdA <= 8'b00110100;
8'b00110101: rdA <= 8'b00110101;
8'b00110110: rdA <= 8'b00110110;
8'b00110111: rdA <= 8'b00110111;
8'b00111000: rdA <= 8'b00111000;
8'b00111001: rdA <= 8'b00111001;
8'b00111010: rdA <= 8'b00111010;
8'b00111011: rdA <= 8'b00111011;
8'b00111100: rdA <= 8'b00111100;
8'b00111101: rdA <= 8'b00111101;
8'b00111110: rdA <= 8'b00111110;
8'b00111111: rdA <= 8'b00111111;
8'b01000000: rdA <= 8'b01000000;
8'b01000001: rdA <= 8'b01000001;
8'b01000010: rdA <= 8'b01000010;
8'b01000011: rdA <= 8'b01000011;
8'b01000100: rdA <= 8'b01000100;
8'b01000101: rdA <= 8'b01000101;
8'b01000110: rdA <= 8'b01000110;
8'b01000111: rdA <= 8'b01000111;
8'b01001000: rdA <= 8'b01001000;
8'b01001001: rdA <= 8'b01001001;
8'b01001010: rdA <= 8'b01001010;
8'b01001011: rdA <= 8'b01001011;
8'b01001100: rdA <= 8'b01001100;
8'b01001101: rdA <= 8'b01001101;
8'b01001110: rdA <= 8'b01001110;
8'b01001111: rdA <= 8'b01001111;
8'b01010000: rdA <= 8'b01010000;
8'b01010001: rdA <= 8'b01010001;
8'b01010010: rdA <= 8'b01010010;
8'b01010011: rdA <= 8'b01010011;
8'b01010100: rdA <= 8'b01010100;
8'b01010101: rdA <= 8'b01010101;
8'b01010110: rdA <= 8'b01010110;
8'b01010111: rdA <= 8'b01010111;
8'b01011000: rdA <= 8'b01011000;
8'b01011001: rdA <= 8'b01011001;
8'b01011010: rdA <= 8'b01011010;
8'b01011011: rdA <= 8'b01011011;
8'b01011100: rdA <= 8'b01011100;
8'b01011101: rdA <= 8'b01011101;
8'b01011110: rdA <= 8'b01011110;
8'b01011111: rdA <= 8'b01011111;
8'b01100000: rdA <= 8'b01100000;
8'b01100001: rdA <= 8'b01100001;
8'b01100010: rdA <= 8'b01100010;
8'b01100011: rdA <= 8'b01100011;
8'b01100100: rdA <= 8'b01100100;
8'b01100101: rdA <= 8'b01100101;
8'b01100110: rdA <= 8'b01100110;
8'b01100111: rdA <= 8'b01100111;
8'b01101000: rdA <= 8'b01101000;
8'b01101001: rdA <= 8'b01101001;
8'b01101010: rdA <= 8'b01101010;
8'b01101011: rdA <= 8'b01101011;
8'b01101100: rdA <= 8'b01101100;
8'b01101101: rdA <= 8'b01101101;
8'b01101110: rdA <= 8'b01101110;
8'b01101111: rdA <= 8'b01101111;
8'b01110000: rdA <= 8'b01110000;
8'b01110001: rdA <= 8'b01110001;
8'b01110010: rdA <= 8'b01110010;
8'b01110011: rdA <= 8'b01110011;
8'b01110100: rdA <= 8'b01110100;
8'b01110101: rdA <= 8'b01110101;
8'b01110110: rdA <= 8'b01110110;
8'b01110111: rdA <= 8'b01110111;
8'b01111000: rdA <= 8'b01111000;
8'b01111001: rdA <= 8'b01111001;
8'b01111010: rdA <= 8'b01111010;
8'b01111011: rdA <= 8'b01111011;
8'b01111100: rdA <= 8'b01111100;
8'b01111101: rdA <= 8'b01111101;
8'b01111110: rdA <= 8'b01111110;
8'b01111111: rdA <= 8'b01111111;
8'b10000000 : rdA <= 8'b10000000;
8'b10000001 : rdA <= 8'b10000001;
8'b10000010 : rdA <= 8'b10000010;
8'b10000011 : rdA <= 8'b10000011;
8'b10000100 : rdA <= 8'b10000100;
8'b10000101 : rdA <= 8'b10000101;
8'b10000110 : rdA <= 8'b10000110;
8'b10000111 : rdA <= 8'b10000111;
8'b10001000 : rdA <= 8'b10001000;
8'b10001001 : rdA <= 8'b10001001;
8'b10001010 : rdA <= 8'b10001010;
8'b10001011 : rdA <= 8'b10001011;
8'b10001100 : rdA <= 8'b10001100;
8'b10001101 : rdA <= 8'b10001101;
8'b10001110 : rdA <= 8'b10001110;
8'b10001111 : rdA <= 8'b10001111;
8'b10010000 : rdA <= 8'b10010000;
8'b10010001 : rdA <= 8'b10010001;
8'b10010010 : rdA <= 8'b10010010;
8'b10010011 : rdA <= 8'b10010011;
8'b10010100 : rdA <= 8'b10010100;
8'b10010101 : rdA <= 8'b10010101;
8'b10010110 : rdA <= 8'b10010110;
8'b10010111 : rdA <= 8'b10010111;
8'b10011000 : rdA <= 8'b10011000;
8'b10011001 : rdA <= 8'b10011001;
8'b10011010 : rdA <= 8'b10011010;
8'b10011011 : rdA <= 8'b10011011;
8'b10011100 : rdA <= 8'b10011100;
8'b10011101 : rdA <= 8'b10011101;
8'b10011110 : rdA <= 8'b10011110;
8'b10011111 : rdA <= 8'b10011111;
8'b10100000 : rdA <= 8'b10100000 ;
8'b10100001 : rdA <= 8'b10100001 ;
8'b10100010 : rdA <= 8'b10100010 ;
8'b10100011 : rdA <= 8'b10100011 ;
8'b10100100 : rdA <= 8'b10100100 ;
8'b10100101 : rdA <= 8'b10100101 ;
8'b10100110 : rdA <= 8'b10100110 ;
8'b10100111 : rdA <= 8'b10100111 ;
8'b10101000 : rdA <= 8'b10101000 ;
8'b10101001 : rdA <= 8'b10101001 ;
8'b10101010 : rdA <= 8'b10101010 ;
8'b10101011 : rdA <= 8'b10101011 ;
8'b10101100 : rdA <= 8'b10101100 ;
8'b10101101 : rdA <= 8'b10101101 ;
8'b10101110 : rdA <= 8'b10101110 ;
8'b10101111 : rdA <= 8'b10101111 ;
8'b10110000 : rdA <= 8'b10110000;
8'b10110001 : rdA <= 8'b10110001;
8'b10110010 : rdA <= 8'b10110010;
8'b10110011 : rdA <= 8'b10110011;
8'b10110100 : rdA <= 8'b10110100;
8'b10110101 : rdA <= 8'b10110101;
8'b10110110 : rdA <= 8'b10110110;
8'b10110111 : rdA <= 8'b10110111;
8'b10111000 : rdA <= 8'b10111000;
8'b10111001 : rdA <= 8'b10111001;
8'b10111010 : rdA <= 8'b10111010;
8'b10111011 : rdA <= 8'b10111011;
8'b10111100 : rdA <= 8'b10111100;
8'b10111101 : rdA <= 8'b10111101;
8'b10111110 : rdA <= 8'b10111110;
8'b10111111 : rdA <= 8'b10111111;
8'b11000000 : rdA <= 8'b11000000;
8'b11000001 : rdA <= 8'b11000001;
8'b11000010 : rdA <= 8'b11000010;
8'b11000011 : rdA <= 8'b11000011;
8'b11000100 : rdA <= 8'b11000100;
8'b11000101 : rdA <= 8'b11000101;
8'b11000110 : rdA <= 8'b11000110;
8'b11000111 : rdA <= 8'b11000111;
8'b11001000 : rdA <= 8'b11001000;
8'b11001001 : rdA <= 8'b11001001;
8'b11001010 : rdA <= 8'b11001010;
8'b11001011 : rdA <= 8'b11001011;
8'b11001100 : rdA <= 8'b11001100;
8'b11001101 : rdA <= 8'b11001101;
8'b11001110 : rdA <= 8'b11001110;
8'b11001111 : rdA <= 8'b11001111;
8'b11010000 : rdA <= 8'b11010000;
8'b11010001 : rdA <= 8'b11010001;
8'b11010010 : rdA <= 8'b11010010;
8'b11010011 : rdA <= 8'b11010011;
8'b11010100 : rdA <= 8'b11010100;
8'b11010101 : rdA <= 8'b11010101;
8'b11010110 : rdA <= 8'b11010110;
8'b11010111 : rdA <= 8'b11010111;
8'b11011000 : rdA <= 8'b11011000;
8'b11011001 : rdA <= 8'b11011001;
8'b11011010 : rdA <= 8'b11011010;
8'b11011011 : rdA <= 8'b11011011;
8'b11011100 : rdA <= 8'b11011100;
8'b11011101 : rdA <= 8'b11011101;
8'b11011110 : rdA <= 8'b11011110;
8'b11011111 : rdA <= 8'b11011111;
8'b11100000 : rdA <= 8'b11100000; 
8'b11100001 : rdA <= 8'b11100001;
8'b11100010 : rdA <= 8'b11100010;
8'b11100011 : rdA <= 8'b11100011;
8'b11100100 : rdA <= 8'b11100100;
8'b11100101 : rdA <= 8'b11100101;
8'b11100110 : rdA <= 8'b11100110;
8'b11100111 : rdA <= 8'b11100111;
8'b11101000 : rdA <= 8'b11101000;
8'b11101001 : rdA <= 8'b11101001;
8'b11101010 : rdA <= 8'b11101010;
8'b11101011 : rdA <= 8'b11101011;
8'b11101100 : rdA <= 8'b11101100;
8'b11101101 : rdA <= 8'b11101101;
8'b11101110 : rdA <= 8'b11101110;
8'b11101111 : rdA <= 8'b11101111;
8'b11110000 : rdA <= 8'b11110000;
8'b11110001 : rdA <= 8'b11110001;
8'b11110010 : rdA <= 8'b11110010;
8'b11110011 : rdA <= 8'b11110011;
8'b11110100 : rdA <= 8'b11110100;
8'b11110101 : rdA <= 8'b11110101;
8'b11110110 : rdA <= 8'b11110110;
8'b11110111 : rdA <= 8'b11110111;
8'b11111000 : rdA <= 8'b11111000;
8'b11111001 : rdA <= 8'b11111001;
8'b11111010 : rdA <= 8'b11111010;
8'b11111011 : rdA <= 8'b11111011;
8'b11111100 : rdA <= 8'b11111100;
8'b11111101 : rdA <= 8'b11111101;
8'b11111110 : rdA <= 8'b11111110;
8'b11111111 : rdA <= 8'b11111111;
endcase
end

always@(posedge clk) begin
rdB <= rdB + 1'b1;
if(rdB > 8'b11111111) begin
  rdB <= 8'b00000000;
end
end
endmodule

module mux_rdA(
input [7:0] rdA,
output reg [7:0] result_rdA
);
reg select_mux;
always@(select_mux) begin
case(select_mux) 
1'b0 : result_rdA <= rdA;
1'b1 : begin result_rdA <= rdA + 1'b1;
if(result_rdA > 8'b11111111) begin
result_rdA <= 8'b00000000;
end
end

endcase
end
endmodule

module mux_rdB(
input [7:0] rdB,
output reg [7:0] result_rdB
);
reg select_mux;
always@(select_mux) begin
case(select_mux) 
1'b0 : result_rdB <= rdB;
1'b1 : begin result_rdB <= rdB + 1'b1;
if(result_rdB > 8'b11111111) begin
result_rdB <= 8'b00000000;
end
end

endcase
end
endmodule
